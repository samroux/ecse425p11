
entity rtl_BLOCKNAME is
   port (
		

   );
end entity rtl_BLOCKNAME;

architecture rtl of rtl_BLOCKNAME is

begin

end architecture rtl;